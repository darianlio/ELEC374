module MDR (clk, clear,